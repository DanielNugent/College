--Daniel Nugent
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY control_memory IS
    PORT (

        IN_CAR : IN std_logic_vector(7 DOWNTO 0);
        MW : OUT std_logic;

        MM : OUT std_logic;

        RW : OUT std_logic;

        MD : OUT std_logic;

        FS : OUT std_logic_vector(4 DOWNTO 0);

        MB : OUT std_logic;

        TB : OUT std_logic;

        TA : OUT std_logic;

        TD : OUT std_logic;

        PL : OUT std_logic;

        PI : OUT std_logic;

        IL : OUT std_logic;

        MC : OUT std_logic;

        MS : OUT std_logic_vector(2 DOWNTO 0);

        NA : OUT std_logic_vector(7 DOWNTO 0)

    );
END control_memory;

ARCHITECTURE Behavioral OF control_memory IS

    TYPE mem_array IS ARRAY(0 TO 255) OF std_logic_vector(27 DOWNTO 0);

BEGIN
    memory_m : PROCESS (IN_CAR)
        VARIABLE control_mem : mem_array := (

        x"C020306",
        x"C02400E",
        x"C020184",
        X"C020054",
        X"0000000",
        X"0000000",
        X"0000000",
        X"0000000",
        X"0000000",
        X"0000000",
        X"0000000",
        X"0000000",
        X"0000000",
        X"0000000",
        X"0000000",
        X"0000000",

        -- Module 1
        X"C030024", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000",

        -- Module 2
        X"0000000", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000",

        -- Module 3
        X"0000000", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000",

        -- Module 4
        X"0000000", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000",

        -- Module 5
        X"0000000", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000",

        -- Module 6
        X"0000000", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000",

        -- Module 7
        X"0000000", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000",

        --  Module 8
        X"0000000", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000",

        -- Module 9
        X"0000000", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000",

        -- Module A
        X"0000000", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000",

        -- Module B
        X"0000000", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000",

        -- Module C
        x"C12C002",
        x"0030000",
        X"0000000",
        X"0000000",
        X"0000000",
        X"0000000",
        X"0000000",
        X"0000000",
        X"0000000",
        X"0000000",
        X"0000000",
        X"0000000",
        X"0000000",
        X"0000000",
        X"0000000",
        X"0000000",

        -- Module D
        X"C10C002",
        X"0030004",
        X"0000000",
        X"0000000",
        X"0000000",
        X"0000000",
        X"0000000",
        X"0000000",
        X"0000000",
        X"0000000",
        X"0000000",
        X"0000000",
        X"0000000",
        X"0000000",
        X"0000000",
        X"0000000",

        -- Module E
        X"0000000", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000",

        -- Module F
        X"0000000", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000",
        X"0000000", X"0000000", X"0000000", X"0000000");

        VARIABLE addr : INTEGER;
        VARIABLE control_out : std_logic_vector(27 DOWNTO 0);

    BEGIN
        addr := conv_integer(IN_CAR);
        control_out := control_mem(addr);

        MW <= control_out(0);
        MM <= control_out(1);
        RW <= control_out(2);
        MD <= control_out(3);
        FS <= control_out(8 DOWNTO 4);
        MB <= control_out(9);
        TB <= control_out(10);
        TA <= control_out(11);
        TD <= control_out(12);
        PL <= control_out(13);
        PI <= control_out(14);
        IL <= control_out(15);
        MC <= control_out(16);
        MS <= control_out(19 DOWNTO 17);
        NA <= control_out(27 DOWNTO 20);
    END PROCESS;

END Behavioral;